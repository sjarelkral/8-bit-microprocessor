`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    19:32:41 06/05/2020
// Design Name:
// Module Name:    Microprocessor
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Microprocessor(
    output clock,
    output [7:0]instruction_address,
    output [6:0]high_reg_write_data,
    output [6:0]low_reg_write_data,
    input oscillator,
    input reset,
    input [7:0]instruction
    );

    //Frequency divider : Generate 1 Hz clock (output LED, internal input for components)
    reg [25:0] delay;
    reg sec;
    always @(posedge oscillator)begin
    	delay  <= (delay == 25000000)?26'd0:(delay+1);
    	if (delay == 26'd0)begin
    		sec <= ~sec;
    	end
    end
    assign clock = sec;

    //Storage elements
    reg [7:0]registers[3:0];
    reg [7:0]pc;
    reg [7:0]ir;
    reg [7:0]memory[31:0];


    always @ (posedge reset or posedge clock) begin

    if (reset) begin
      //reset pc
      pc <= 8'd0;

      //reset registers
      registers <= 32'd0;

      //reinitialize memory
      memory[0] <= 8'd0;
      memory[1] <= 8'd1;
      memory[2] <= 8'd2;
      memory[3] <= 8'd3;
      memory[4] <= 8'd4;
      memory[5] <= 8'd5;
      memory[6] <= 8'd6;
      memory[7] <= 8'd7;
      memory[8] <= 8'd8;
      memory[9] <= 8'd9;
      memory[10] <= 8'd10;
      memory[11] <= 8'd11;
      memory[12] <= 8'd12;
      memory[13] <= 8'd13;
      memory[14] <= 8'd14;
      memory[15] <= 8'd15;
      memory[16] <= 8'd0;
      memory[17] <= 8'd-1;
      memory[18] <= 8'd-2;
      memory[19] <= 8'd-3;
      memory[20] <= 8'd-4;
      memory[21] <= 8'd-5;
      memory[22] <= 8'd-6;
      memory[23] <= 8'd-7;
      memory[24] <= 8'd-8;
      memory[25] <= 8'd-9;
      memory[26] <= 8'd-10;
      memory[27] <= 8'd-11;
      memory[28] <= 8'd-12;
      memory[29] <= 8'd-13;
      memory[30] <= 8'd-14;
      memory[31] <= 8'd-15;
    end


    end











    reg [7:0]console_buffer;

    Console disp1(high_out, console_buffer[7:4]);
    Console disp2(low_out, console_buffer[3:0]);

	 //Buses
	 wire RegDst;
   wire RegWrite;
   wire ALUSrc;
   wire Branch;
   wire MemRead;
   wire MemWrite;
   wire MemtoReg;
   wire ALUOp;
   wire [1:0]ReadRegister1;
   wire [1:0]ReadRegister2;
   wire [1:0]WriteRegister;
	 wire [7:0]MemAddress;
   wire [7:0]ALUResult;
   wire [7:0]ALUin1;
   wire [7:0]ALUin2;
	 wire [7:0]ReadData1; //reg
	 wire [7:0]ReadData2; //reg
	 wire [7:0]ReadData; //mem
	 wire [7:0]RegWriteData;
	 wire [7:0]WriteData;
	 wire [7:0]SignExtImm;





   //PC
   assign PCAddess = PC; // Instruction  = Instruction Memory[PC]

   //Instruction OP code is used to generate control signals
   assign RegDst =  ~IR[6];
	 assign RegWrite = ~IR[7];
	 assign ALUSrc = IR[7] ^ IR[6];
	 assign Branch  = IR[7]& IR[6];
	 assign MemRead = (IR[7:6] == 2'b01 );
	 assign MemWrite = (IR[7:6] == 2'b10);
	 assign MemtoReg = IR[6];
	 assign ALUOp = ~(IR[7] | IR[6]);

   //Register input/output connections
   assign ReadRegister1 = IR[5:4];
   assign ReadRegister2 = IR[3:2];
   assign WriteRegister = RegDst ? IR[1:0] : IR[3:2];
   assign RegWriteData = (MemtoReg) ? ReadData : ALUResult;

   assign ReadData1 = (ReadRegister1 == 2'd0) ? GPR[0]:
                      (ReadRegister1 == 2'd1) ? GPR[1]:
                      (ReadRegister1 == 2'd2) ? GPR[2]:
							 GPR[3];

    assign ReadData2 = (ReadRegister2 == 2'd0) ? GPR[0]:
                      (ReadRegister2 == 2'd1) ? GPR[1]:
                      (ReadRegister2 == 2'd2) ? GPR[2]:
							 GPR[3];


   //Sign extend Instruction [1:0]
   assign SignExtImm[1:0] = IR[1:0];
   assign SignExtImm[7:2] = (IR[1]) ? 6'b111111 : 6'b000000;

   //connections into the ALU
   assign ALUin1  = ReadData1;
   assign ALUin2 = (ALUSrc) ? SignExtImm : ReadData2;
   assign ALUResult = ALUin1 + ALUin2;

   //Memory input/output values
   assign MemAddress = ALUResult;
   assign WriteData = ReadData2;
   assign ReadData = DataMemory[MemAddress];

   always @ ( posedge clock or posedge reset) begin
      if (reset)begin

        //Reset PC
        PC <= 8'd0;

        //Reset registers
        GPR[0] <= 8'd0;
        GPR[1] <= 8'd0;
        GPR[2] <= 8'd0;
        GPR[3] <= 8'd0;

         //Reinitialize memory;
         DataMemory[0] <= 8'd0;
         DataMemory[1] <= 8'd1;
         DataMemory[2] <= 8'd2;
         DataMemory[3] <= 8'd3;
         DataMemory[4] <= 8'd4;
         DataMemory[5] <= 8'd5;
         DataMemory[6] <= 8'd6;
         DataMemory[7] <= 8'd7;
         DataMemory[8] <= 8'd8;
         DataMemory[9] <= 8'd9;
         DataMemory[10] <= 8'd10;
         DataMemory[11] <= 8'd11;
         DataMemory[12] <= 8'd12;
         DataMemory[13] <= 8'd13;
         DataMemory[14] <= 8'd14;
         DataMemory[15] <= 8'd15;
         DataMemory[16] <= 8'd16;
         DataMemory[17] <= 8'd17;
         DataMemory[18] <= 8'd18;
         DataMemory[19] <= 8'd19;
         DataMemory[20] <= 8'd20;
         DataMemory[21] <= 8'd21;
         DataMemory[22] <= 8'd22;
         DataMemory[23] <= 8'd23;
         DataMemory[24] <= 8'd24;
         DataMemory[25] <= 8'd25;
         DataMemory[26] <= 8'd26;
         DataMemory[27] <= 8'd27;
         DataMemory[28] <= 8'd28;
         DataMemory[29] <= 8'd29;
         DataMemory[30] <= 8'd30;
         DataMemory[31] <= 8'd31;
       end

       else begin

       IR <= Instruction;
       PC <= Branch ? PC+1+SignExtImm : PC+1; //Evaluate PC

       if (RegWrite) begin
         case (WriteRegister)
           2'd0: GPR[0] <= RegWriteData;
           2'd1: GPR[1] <= RegWriteData;
           2'd2: GPR[2] <= RegWriteData;
           2'd3: GPR[3] <= RegWriteData;
         endcase
         console_buffer <= RegWriteData;
       end

       if (MemWrite) begin
         DataMemory[MemAddress] <= WriteData;
       end
		 end

		 end

endmodule
